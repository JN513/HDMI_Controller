module top (
    input  logic clk,
    input  logic rst_i,

    output logic TXD,
    input  logic RXD,

    output logic [5:0]led
);




endmodule
